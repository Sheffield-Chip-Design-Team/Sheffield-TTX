/*
 * Copyright (c) 2024 - James Ashie Kotey
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

// BUILD TIME: 2024-11-30 19:42:10.694939 

module tt_um_vga_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

//using full adder
  FullAdder fa (.a(ui_in[0]), .b(ui_in[1]), .c(ui_in[2]), .carry(uo_out[1]), .sum(uo_out[0]));

  // All output pins must be assigned. If not used, assign to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;
  assign uo_out[7:2] = 0;
    
endmodule

//================================================
//Module: Full Adder Verilog Code
//Author(s): James Ashie Kotey 
//Last Updated:  8/5/24

module FullAdder(a,b,c, sum, carry);
    
    //Ports
    input a,b,c;
    output sum,carry;
    
    //Implimentation
    assign sum = (a^b)^ c;
    assign carry = (((a^b)&c) | (a&b)); // Use | for Or Not +

endmodule

