// Game control Unit
// Last Updated: 31/01/2025 @ 16:23:52

module GameStateControlUnit (
    input             clk,
    input wire [7:0]  playerPos,
    input wire [55:0] dragonSegmentPositions

);






endmodule