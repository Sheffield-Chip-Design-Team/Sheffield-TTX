// Game control Unit
// Last Updated: 

module GameStateControlUnit (
    input             clk,
    input wire [7:0]  playerPos,
    input wire [55:0] dragonSegmentPositions

);






endmodule