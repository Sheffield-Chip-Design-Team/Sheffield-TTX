
// Module : Sheep Logic

// coordinate system  
// location [7:0]
// location [7:4] - the x coordinates
// location [3:0] - the y coordinates
// the limits for the screen are (0,0) - > (15,11)

module sheepLogic (
    input clk,
    input reset,
    input wire read_enable, // When high, generate random position for the sheep
    input wire [7:0] dragon_pos, // using as seed value to ensure no overlap
    input wire [7:0] player_pos, // using as seed value to ensure no overlap
    output reg [7:0] sheep_pos, // 8-bit position (4 bits for X, 4 bits for Y)
    output reg [3:0] sheep_sprite
);

    wire [7:0] random_value; // 8-bit random value: first 4 bits -> X, last 4 bits -> Y

    // Instantiate the random number generator with seeded initial value
    rand_num rng (
        .clk(clk),
        .reset(reset),
        .seed((player_pos ^ dragon_pos) + 1'b1), // Seed with XOR of player and dragon positions +1
        .rdm_num(random_value)                // Random value generated by the RNG

    );

    always @(posedge clk) begin
        if (~reset) begin
        
            if (read_enable) begin
                sheep_sprite <= 1; 
                // Generate a valid position
                // add masks to enforce limit
                sheep_pos[7:4] <= random_value[7:4];

                // enforce limit 
                if (random_value[3:0] > 11) begin // can probably be minimised
                    sheep_pos[3:0] <= ~random_value[3:0];
                end else begin
                    sheep_pos[3:0] <= random_value[3:0];
                end
            end
        
        end else begin
            // Reset condition: sheep is not visible and position off-screen
            sheep_sprite <= 0;
            // sheep_pos <= 8'b0; // Initialize to 0 during reset
        end
    end
    /*

        y position  correction
            0000       - 
            0001       -
            0010       -
            0011       -
            0100       -
            0101       -
            0110       -
            0111       -
            1000       -
            1001       -
            1010       -
            1011       -
            1100       0011
            1101       0010
            1110       0001  
            1111       0000
    */

    endmodule

    module rand_num (
        input wire clk,
        input wire reset,
        input wire [7:0] seed, // Seed input for initializing randomness
        output reg [7:0] rdm_num
    );

    reg [2:0] counter;

    always @(posedge clk or posedge reset) begin
        
        if (reset) begin // for when we need a new random immediately
            rdm_num <= seed;  // Initialize value using the trigger
            counter <= 7;     // Reset counter
        
        end else if (counter > 0) begin
            // Shift and apply feedback for randomness
            rdm_num[6:0] <= rdm_num[7:1];  // Shift all bits
            rdm_num[7] <= rdm_num[6] ^ rdm_num[5] ^ rdm_num[4]; // Feedback XOR for randomness
            counter <= counter - 1;        // Decrement counter

        end else begin
            counter <= 7;  // Reset counter for next random number
            rdm_num <= seed;
        end
    end

endmodule



